library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity temporizador is
    generic (
        N : integer);
    port (
        clk : in std_logic;
        hab : in std_logic;
        reset : in std_logic;
        reset_emergencia: in std_logic;

        P : in std_logic_vector (N-1 downto 0);
        Z : out std_logic;
        T : out std_logic);
end temporizador;

architecture arch of temporizador is
    signal D, D_sig : unsigned (N-1 downto 0);
begin

    memoria : process (clk)
    begin
        if rising_edge(clk) then
            D <= D_sig;
        end if;
    end process;

    D_sig <= to_unsigned(1, N) when reset_emergencia else
            (others=>'0') when reset else
             D when not hab else
             unsigned(P) when Z else
             D - 1;
    Z <= D ?= 0;
    T <= D ?= 1;
end arch;
